configuration xor_conf of XOR_GATE is

    for behaviour
    end for;

end;
