package t is end;

package body t is

    procedure t is
    begin
	while TRUE loop
	    exit when FALSE;
	end loop;
    end;

end;
