architecture hallo of huhu is
begin
end;
