entity huhu is
end;
