--*- text -*-

package beispiel is

    function main ( signal x: integer ) return integer;

    constant pi : real;

end;
