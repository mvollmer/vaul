configuration anderer_half_adder of half_adder is

    for structure
	for all : AND_GATE
    	    generic map ( 100 ns );
	end for;
    end for;

end;
